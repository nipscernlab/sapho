module rel_addr
#(
	parameter MDATAW = 8,
	parameter FFTSIZ = 3,

	parameter USEFFT = 1
)
(
	input               srf, inv,
	input  [MDATAW-1:0] in,
	input  [MDATAW-1:0] addr,
	output [MDATAW-1:0] out
);

generate 

	if (USEFFT) begin

		reg [FFTSIZ-1:0] aux;

		integer i;

		always @ (*) begin
			for (i = 0; i < FFTSIZ; i = i+1) begin : norm
				aux[i] <= in[FFTSIZ-i];
			end
		end

		//pula o LSB para pegar real e imaginario em sequencia
		wire [MDATAW-1:0] add = (inv) ? {in[MDATAW-1:FFTSIZ+1], aux, in[0]} : in;

		assign out = (srf) ? add + addr: addr;

	end else

		assign out = (srf) ? in  + addr: addr;

endgenerate

endmodule 